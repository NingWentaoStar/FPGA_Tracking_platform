module median_filter(

   );
endmodule